module lol-qwop ;
   
  initial begin
    $display ("lol-qwop");
    $finish;
  end
  
endmodule 
